module mux_16X1_32bit(
		input  logic [3:0] sel,
		input  logic [31:0] D0, D1, D2, D3, D4, D5, D6, D7, D8,
        input  logic [31:0] D9, D10, D11, D12, D13, D14, D15,
		output logic [31:0] Y
);

//This is an intientional error: the 8-bit input D is writen in reversed this whole time
//Consider modify the module that already adapt to the previous issued version



mux_16X1   bit0(.sel(sel), .Y(Y[0]),   .D({D15[0], D14[0], D13[0],  D12[0],  D11[0],  D10[0],  D9[0],  D8[0],
                                           D7[0],  D6[0],  D5[0],   D4[0],   D3[0],   D2[0],   D1[0],  D0[0]}));
															
mux_16X1   bit1(.sel(sel), .Y(Y[1]),   .D({D15[1], D14[1], D13[1],  D12[1],  D11[1],  D10[1],  D9[1],  D8[1],
                                           D7[1],  D6[1],  D5[1],   D4[1],   D3[1],   D2[1],   D1[1],  D0[1]}));

mux_16X1   bit2(.sel(sel), .Y(Y[2]),   .D({D15[2], D14[2], D13[2],  D12[2],  D11[2],  D10[2],  D9[2],  D8[2],
                                           D7[2],  D6[2],  D5[2],   D4[2],   D3[2],   D2[2],   D1[2],  D0[2]}));

mux_16X1   bit3(.sel(sel), .Y(Y[3]),   .D({D15[3], D14[3], D13[3],  D12[3],  D11[3],  D10[3],  D9[3],  D8[3],
                                           D7[3],  D6[3],  D5[3],   D4[3],   D3[3],   D2[3],   D1[3],  D0[3]}));

mux_16X1   bit4(.sel(sel), .Y(Y[4]),   .D({D15[4], D14[4], D13[4],  D12[4],  D11[4],  D10[4],  D9[4],  D8[4],
                                           D7[4],  D6[4],  D5[4],   D4[4],   D3[4],   D2[4],   D1[4],  D0[4]}));

mux_16X1   bit5(.sel(sel), .Y(Y[5]),   .D({D15[5], D14[5], D13[5],  D12[5],  D11[5],  D10[5],  D9[5],  D8[5],
                                           D7[5],  D6[5],  D5[5],   D4[5],   D3[5],   D2[5],   D1[5],  D0[5]}));
															
mux_16X1   bit6(.sel(sel), .Y(Y[6]),   .D({D15[6], D14[6], D13[6],  D12[6],  D11[6],  D10[6],  D9[6],  D8[6],
                                           D7[6],  D6[6],  D5[6],   D4[6],   D3[6],   D2[6],   D1[6],  D0[6]}));
															
mux_16X1   bit7(.sel(sel), .Y(Y[7]),   .D({D15[7], D14[7], D13[7],  D12[7],  D11[7],  D10[7],  D9[7],  D8[7],
                                           D7[7],  D6[7],  D5[7],   D4[7],   D3[7],   D2[7],   D1[7],  D0[7]}));
															
mux_16X1   bit8(.sel(sel), .Y(Y[8]),   .D({D15[8], D14[8], D13[8],  D12[8],  D11[8],  D10[8],  D9[8],  D8[8],
                                           D7[8],  D6[8],  D5[8],   D4[8],   D3[8],   D2[8],   D1[8],  D0[8]}));
															
mux_16X1   bit9(.sel(sel), .Y(Y[9]),   .D({D15[9], D14[9], D13[9],  D12[9],  D11[9],  D10[9],  D9[9],  D8[9],
                                           D7[9],  D6[9],  D5[9],   D4[9],   D3[9],   D2[9],   D1[9],  D0[9]}));
															
mux_16X1   bit10(.sel(sel), .Y(Y[10]), .D({D15[10], D14[10], D13[10],  D12[10],  D11[10],  D10[10],  D9[10],  D8[10],
                                           D7[10],  D6[10],  D5[10],   D4[10],   D3[10],   D2[10],   D1[10],  D0[10]}));
															 
mux_16X1   bit11(.sel(sel), .Y(Y[11]), .D({D15[11], D14[11], D13[11],  D12[11],  D11[11],  D10[11],  D9[11],  D8[11],
                                           D7[11],  D6[11],  D5[11],   D4[11],   D3[11],   D2[11],   D1[11],  D0[11]}));
															 
mux_16X1   bit12(.sel(sel), .Y(Y[12]), .D({D15[12], D14[12], D13[12],  D12[12],  D11[12],  D10[12],  D9[12],  D8[12],
                                           D7[12],  D6[12],  D5[12],   D4[12],   D3[12],   D2[12],   D1[12],  D0[12]}));
															 
mux_16X1   bit13(.sel(sel), .Y(Y[13]), .D({D15[13], D14[13], D13[13],  D12[13],  D11[13],  D10[13],  D9[13],  D8[13],
                                           D7[13],  D6[13],  D5[13],   D4[13],   D3[13],   D2[13],   D1[13],  D0[13]}));
															 
mux_16X1   bit14(.sel(sel), .Y(Y[14]), .D({D15[14], D14[14], D13[14],  D12[14],  D11[14],  D10[14],  D9[14],  D8[14],
                                           D7[14],  D6[14],  D5[14],   D4[14],   D3[14],   D2[14],   D1[14],  D0[14]}));
															 
mux_16X1   bit15(.sel(sel), .Y(Y[15]), .D({D15[15], D14[15], D13[15],  D12[15],  D11[15],  D10[15],  D9[15],  D8[15],
                                           D7[15],  D6[15],  D5[15],   D4[15],   D3[15],   D2[15],   D1[15],  D0[15]}));
															  
mux_16X1   bit16(.sel(sel), .Y(Y[16]), .D({D15[16], D14[16], D13[16],  D12[16],  D11[16],  D10[16],  D9[16],  D8[16],
                                           D7[16],  D6[16],  D5[16],   D4[16],   D3[16],   D2[16],   D1[16],  D0[16]}));
															  
mux_16X1   bit17(.sel(sel), .Y(Y[17]), .D({D15[17], D14[17], D13[17],  D12[17],  D11[17],  D10[17],  D9[17],  D8[17],
                                           D7[17],  D6[17],  D5[17],   D4[17],   D3[17],   D2[17],   D1[17],  D0[17]}));
															  
mux_16X1   bit18(.sel(sel), .Y(Y[18]), .D({D15[18], D14[18], D13[18],  D12[18],  D11[18],  D10[18],  D9[18],  D8[18],
                                           D7[18],  D6[18],  D5[18],   D4[18],   D3[18],   D2[18],   D1[18],  D0[18]}));
															  
mux_16X1   bit19(.sel(sel), .Y(Y[19]), .D({D15[19], D14[19], D13[19],  D12[19],  D11[19],  D10[19],  D9[19],  D8[19],
                                           D7[19],  D6[19],  D5[19],   D4[19],   D3[19],   D2[19],   D1[19],  D0[19]}));
															  
mux_16X1   bit20(.sel(sel), .Y(Y[20]), .D({D15[20], D14[20], D13[20],  D12[20],  D11[20],  D10[20],  D9[20],  D8[20],
                                           D7[20],  D6[20],  D5[20],   D4[20],   D3[20],   D2[20],   D1[20],  D0[20]}));
															 
mux_16X1   bit21(.sel(sel), .Y(Y[21]), .D({D15[21], D14[21], D13[21],  D12[21],  D11[21],  D10[21],  D9[21],  D8[21],
                                           D7[21],  D6[21],  D5[21],   D4[21],   D3[21],   D2[21],   D1[21],  D0[21]}));
															 
mux_16X1   bit22(.sel(sel), .Y(Y[22]), .D({D15[22], D14[22], D13[22],  D12[22],  D11[22],  D10[22],  D9[22],  D8[22],
                                           D7[22],  D6[22],  D5[22],   D4[22],   D3[22],   D2[22],   D1[22],  D0[22]}));
															 
mux_16X1   bit23(.sel(sel), .Y(Y[23]), .D({D15[23], D14[23], D13[23],  D12[23],  D11[23],  D10[23],  D9[23],  D8[23],
                                           D7[23],  D6[23],  D5[23],   D4[23],   D3[23],   D2[23],   D1[23],  D0[23]}));
															 
mux_16X1   bit24(.sel(sel), .Y(Y[24]), .D({D15[24], D14[24], D13[24],  D12[24],  D11[24],  D10[24],  D9[24],  D8[24],
                                           D7[24],  D6[24],  D5[24],   D4[24],   D3[24],   D2[24],   D1[24],  D0[24]}));
															 
mux_16X1   bit25(.sel(sel), .Y(Y[25]), .D({D15[25], D14[25], D13[25],  D12[25],  D11[25],  D10[25],  D9[25],  D8[25],
                                           D7[25],  D6[25],  D5[25],   D4[25],   D3[25],   D2[25],   D1[25],  D0[25]}));
															 
mux_16X1   bit26(.sel(sel), .Y(Y[26]), .D({D15[26], D14[26], D13[26],  D12[26],  D11[26],  D10[26],  D9[26],  D8[26],
                                           D7[26],  D6[26],  D5[26],   D4[26],   D3[26],   D2[26],   D1[26],  D0[26]}));
															 
mux_16X1   bit27(.sel(sel), .Y(Y[27]), .D({D15[27], D14[27], D13[27],  D12[27],  D11[27],  D10[27],  D9[27],  D8[27],
                                           D7[27],  D6[27],  D5[27],   D4[27],   D3[27],   D2[27],   D1[27],  D0[27]}));
															 
mux_16X1   bit28(.sel(sel), .Y(Y[28]), .D({D15[28], D14[28], D13[28],  D12[28],  D11[28],  D10[28],  D9[28],  D8[28],
                                           D7[28],  D6[28],  D5[28],   D4[28],   D3[28],   D2[28],   D1[28],  D0[28]}));
															 
mux_16X1   bit29(.sel(sel), .Y(Y[29]), .D({D15[29], D14[29], D13[29],  D12[29],  D11[29],  D10[29],  D9[29],  D8[29],
                                           D7[29],  D6[29],  D5[29],   D4[29],   D3[29],   D2[29],   D1[29],  D0[29]}));
															 
mux_16X1   bit30(.sel(sel), .Y(Y[30]), .D({D15[30], D14[30], D13[30],  D12[30],  D11[30],  D10[30],  D9[30],  D8[30],
                                           D7[30],  D6[30],  D5[30],   D4[30],   D3[30],   D2[30],   D1[30],  D0[30]}));
															 
mux_16X1   bit31(.sel(sel), .Y(Y[31]), .D({D15[31], D14[31], D13[31],  D12[31],  D11[31],  D10[31],  D9[31],  D8[31],
                                           D7[31],  D6[31],  D5[31],   D4[31],   D3[31],   D2[31],   D1[31],  D0[31]}));
															 
endmodule

