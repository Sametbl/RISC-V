module demux_1X2(

    	input  logic D,
	input  logic [3:0] sel,
	output logic [15:0] S
);
