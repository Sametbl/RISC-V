module alu(
		input  logic [3:0]  alu_op,			
		input  logic [31:0] operand_a, operand_b,
		output logic [31:0] alu_data
);
wire logic [31:0] ADD_SUB, SLT_U, XOR, OR, AND, Shift, Reserved;
wire logic [1:0] Shift_mode;
wire logic Sub_mode, SLTU_mode;

assign Reserved      = 32'b0;
assign SLT_U[31:1]   = 31'b0;
assign Sub_mode      = ~alu_op[3] & ~alu_op[2] & ~alu_op[1] &  alu_op[0];  // When alu_op == 4'b0001
assign SLTU_mode     = ~alu_op[3] & ~alu_op[2] &  alu_op[1] &  alu_op[0];  // When alu_op == 4'b0011

// mode = 2'b00 : shift Right logic (default) , when alu_op == 4'b1000
// mode = 2;b01 : shift Left  logic           , when alu_op == 4'b0111
// mode = 2'b10 : shift Right Arithmetic      , when alu_op == 4'b1001
// mode = 2'b11 : Reserved
assign Shift_mode[0] = ~alu_op[3] &  alu_op[2] &  alu_op[1] &  alu_op[0]; //(4'b0111)
assign Shift_mode[1] =  alu_op[3] & ~alu_op[2] & ~alu_op[1] &  alu_op[0]; //(4'b1001)

// Datapath
full_adder_32bit  Ins_ADD_SUB (.A(operand_a), .B(operand_b), .Invert_B(Sub_mode),  .C_in(Sub_mode), .Sum(ADD_SUB), .C_out() );
comparator_32bit  Ins_SLT_U   (.A(operand_a), .B(operand_b), .is_unsigned(SLTU_mode), .smaller(SLT_U[0]), .equal(), .larger() );
shifter_32bit     Ins_S_3mode (.data_in(operand_a), .shift_amount(operand_b[4:0]), .mode(Shift_mode), .data_out(Shift) );
assign OR  = operand_a | operand_b;
assign AND = operand_a & operand_b;
assign XOR = operand_a ^ operand_b;


mux_16X1_32bit	  ALU_out     (.sel(alu_op), .Y(alu_data),
                               .D0(ADD_SUB),   .D1(ADD_SUB),   .D2(SLT_U),     .D3(SLT_U),
                               .D4(XOR),       .D5(OR),        .D6(AND),       .D7(Shift),
                               .D8(Shift),     .D9(Shift),     .D10(Reserved), .D11(Reserved),
			      			   .D12(Reserved), .D13(Reserved), .D14(Reserved), .D15(Reserved)	);


endmodule


