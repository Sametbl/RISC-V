module mux_32X1_32bit(
		input  logic [31:0] D0, D1, D2, D3, D4, D5, D6, D7, D8, D9, D10, D11, D12, D13, D14, D15, D16,
		input  logic [31:0] D17, D18, D19, D20, D21, D22, D23, D24, D25, D26, D27, D28, D29, D30, D31,
		input  logic [4:0] sel,
		output logic [31:0] Y
);

mux_32X1   bit0(.sel(sel), .Y(Y[0]), .D({ D31[0], D30[0],  D29[0], D28[0], D27[0], D26[0], D25[0], D24[0],
                                          D23[0], D22[0],  D21[0], D20[0], D19[0], D18[0], D17[0], D16[0],
                                          D15[0], D14[0],  D13[0], D12[0], D11[0], D10[0], D9[0],  D8[0],
                                          D7[0],  D6[0],   D5[0],  D4[0],  D3[0],  D2[0],  D1[0],  D0[0]}));

mux_32X1   bit1(.sel(sel), .Y(Y[1]), .D({ D31[1], D30[1],  D29[1], D28[1], D27[1], D26[1], D25[1], D24[1],
                                          D23[1], D22[1],  D21[1], D20[1], D19[1], D18[1], D17[1], D16[1],
                                          D15[1], D14[1],  D13[1], D12[1], D11[1], D10[1], D9[1],  D8[1],
                                          D7[1],  D6[1],   D5[1],  D4[1],  D3[1],  D2[1],  D1[1],  D0[1]}));

mux_32X1   bit2(.sel(sel), .Y(Y[2]), .D({ D31[2], D30[2],  D29[2], D28[2], D27[2], D26[2], D25[2], D24[2],
                                          D23[2], D22[2],  D21[2], D20[2], D19[2], D18[2], D17[2], D16[2],
                                          D15[2], D14[2],  D13[2], D12[2], D11[2], D10[2], D9[2],  D8[2],
                                          D7[2],  D6[2],   D5[2],  D4[2],  D3[2],  D2[2],  D1[2],  D0[2]}));

mux_32X1   bit3(.sel(sel), .Y(Y[3]), .D({ D31[3], D30[3],  D29[3], D28[3], D27[3], D26[3], D25[3], D24[3],
                                          D23[3], D22[3],  D21[3], D20[3], D19[3], D18[3], D17[3], D16[3],
                                          D15[3], D14[3],  D13[3], D12[3], D11[3], D10[3], D9[3],  D8[3],
                                          D7[3],  D6[3],   D5[3],  D4[3],  D3[3],  D2[3],  D1[3],  D0[3]}));

mux_32X1   bit4(.sel(sel), .Y(Y[4]), .D({ D31[4], D30[4],  D29[4], D28[4], D27[4], D26[4], D25[4], D24[4],
                                          D23[4], D22[4],  D21[4], D20[4], D19[4], D18[4], D17[4], D16[4],
                                          D15[4], D14[4],  D13[4], D12[4], D11[4], D10[4], D9[4],  D8[4],
                                          D7[4],  D6[4],   D5[4],  D4[4],  D3[4],  D2[4],  D1[4],  D0[4]}));

mux_32X1   bit5(.sel(sel), .Y(Y[5]), .D({ D31[5], D30[5],  D29[5], D28[5], D27[5], D26[5], D25[5], D24[5],
                                          D23[5], D22[5],  D21[5], D20[5], D19[5], D18[5], D17[5], D16[5],
                                          D15[5], D14[5],  D13[5], D12[5], D11[5], D10[5], D9[5],  D8[5],
                                          D7[5],  D6[5],   D5[5],  D4[5],  D3[5],  D2[5],  D1[5],  D0[5]}));
															
mux_32X1   bit6(.sel(sel), .Y(Y[6]), .D({ D31[6], D30[6],  D29[6], D28[6], D27[6], D26[6], D25[6], D24[6],
                                          D23[6], D22[6],  D21[6], D20[6], D19[6], D18[6], D17[6], D16[6],
                                          D15[6], D14[6],  D13[6], D12[6], D11[6], D10[6], D9[6],  D8[6],
                                          D7[6],  D6[6],   D5[6],  D4[6],  D3[6],  D2[6],  D1[6],  D0[6]}));
															
mux_32X1   bit7(.sel(sel), .Y(Y[7]), .D({ D31[7], D30[7],  D29[7], D28[7], D27[7], D26[7], D25[7], D24[7],
                                          D23[7], D22[7],  D21[7], D20[7], D19[7], D18[7], D17[7], D16[7],
                                          D15[7], D14[7],  D13[7], D12[7], D11[7], D10[7], D9[7],  D8[7],
                                          D7[7],  D6[7],   D5[7],  D4[7],  D3[7],  D2[7],  D1[7],  D0[7]}));
															
mux_32X1   bit8(.sel(sel), .Y(Y[8]), .D({ D31[8], D30[8],  D29[8], D28[8], D27[8], D26[8], D25[8], D24[8],
                                          D23[8], D22[8],  D21[8], D20[8], D19[8], D18[8], D17[8], D16[8],
                                          D15[8], D14[8],  D13[8], D12[8], D11[8], D10[8], D9[8],  D8[8],
                                          D7[8],  D6[8],   D5[8],  D4[8],  D3[8],  D2[8],  D1[8],  D0[8]}));
															
mux_32X1   bit9(.sel(sel), .Y(Y[9]), .D({ D31[9], D30[9],  D29[9], D28[9], D27[9], D26[9], D25[9], D24[9],
                                          D23[9], D22[9],  D21[9], D20[9], D19[9], D18[9], D17[9], D16[9],
                                          D15[9], D14[9],  D13[9], D12[9], D11[9], D10[9], D9[9],  D8[9],
                                          D7[9],  D6[9],   D5[9],  D4[9],  D3[9],  D2[9],  D1[9],  D0[9]}));
															
mux_32X1   bit10(.sel(sel), .Y(Y[10]), .D({ D31[10], D30[10],  D29[10], D28[10], D27[10], D26[10], D25[10], D24[10],
                                            D23[10], D22[10],  D21[10], D20[10], D19[10], D18[10], D17[10], D16[10],
                                            D15[10], D14[10],  D13[10], D12[10], D11[10], D10[10], D9[10],  D8[10],
                                            D7[10],  D6[10],   D5[10],  D4[10],  D3[10],  D2[10],  D1[10],  D0[10]}));
															 
mux_32X1   bit11(.sel(sel), .Y(Y[11]), .D({ D31[11], D30[11],  D29[11], D28[11], D27[11], D26[11], D25[11], D24[11],
                                            D23[11], D22[11],  D21[11], D20[11], D19[11], D18[11], D17[11], D16[11],
                                            D15[11], D14[11],  D13[11], D12[11], D11[11], D10[11], D9[11],  D8[11],
                                            D7[11],  D6[11],   D5[11],  D4[11],  D3[11],  D2[11],  D1[11],  D0[11]}));
															 
mux_32X1   bit12(.sel(sel), .Y(Y[12]), .D({ D31[12], D30[12],  D29[12], D28[12], D27[12], D26[12], D25[12], D24[12],
                                            D23[12], D22[12],  D21[12], D20[12], D19[12], D18[12], D17[12], D16[12],
                                            D15[12], D14[12],  D13[12], D12[12], D11[12], D10[12], D9[12],  D8[12],
                                            D7[12],  D6[12],   D5[12],  D4[12],  D3[12],  D2[12],  D1[12],  D0[12]}));
															 
mux_32X1   bit13(.sel(sel), .Y(Y[13]), .D({ D31[13], D30[13], D29[13],  D28[13], D27[13], D26[13], D25[13], D24[13],
                                            D23[13], D22[13],   D21[13], D20[13], D19[13], D18[13], D17[13], D16[13],
                                            D15[13], D14[13],  D13[13], D12[13], D11[13], D10[13], D9[13],  D8[13],
                                            D7[13],  D6[13],   D5[13],  D4[13],  D3[13],  D2[13],  D1[13],  D0[13]}));
															 
mux_32X1   bit14(.sel(sel), .Y(Y[14]), .D({ D31[14], D30[14],  D29[14], D28[14], D27[14], D26[14], D25[14], D24[14],
                                            D23[14], D22[14],  D21[14], D20[14], D19[14], D18[14], D17[14], D16[14],
                                            D15[14], D14[14],  D13[14], D12[14], D11[14], D10[14], D9[14],  D8[14],
                                            D7[14],  D6[14],   D5[14],  D4[14],  D3[14],  D2[14],  D1[14],  D0[14]}));
															 
mux_32X1   bit15(.sel(sel), .Y(Y[15]), .D({ D31[15], D30[15],  D29[15], D28[15], D27[15], D26[15], D25[15], D24[15],
                                            D23[15], D22[15],  D21[15], D20[15], D19[15], D18[15], D17[15], D16[15],
                                            D15[15], D14[15],  D13[15], D12[15], D11[15], D10[15], D9[15],  D8[15],
                                            D7[15],  D6[15],   D5[15],  D4[15],  D3[15],  D2[15],  D1[15],  D0[15]}));
															 
mux_32X1   bit16(.sel(sel), .Y(Y[16]), .D({ D31[16], D30[16],  D29[16], D28[16], D27[16], D26[16], D25[16], D24[16],
                                            D23[16], D22[16],  D21[16], D20[16], D19[16], D18[16], D17[16], D16[16],
                                            D15[16], D14[16],  D13[16], D12[16], D11[16], D10[16], D9[16],  D8[16],
                                            D7[16],  D6[16],   D5[16],  D4[16],  D3[16],  D2[16],  D1[16],  D0[16]}));
															 
mux_32X1   bit17(.sel(sel), .Y(Y[17]), .D({ D31[17], D30[17],  D29[17], D28[17], D27[17], D26[17], D25[17], D24[17],
                                            D23[17], D22[17],  D21[17], D20[17], D19[17], D18[17], D17[17], D16[17],
                                            D15[17], D14[17],  D13[17], D12[17], D11[17], D10[17], D9[17],  D8[17],
                                            D7[17],  D6[17],   D5[17],  D4[17],  D3[17],  D2[17],  D1[17],  D0[17]}));
															 
mux_32X1   bit18(.sel(sel), .Y(Y[18]), .D({ D31[18], D30[18],  D29[18], D28[18], D27[18], D26[18], D25[18], D24[18],
                                            D23[18], D22[18],  D21[18], D20[18], D19[18], D18[18], D17[18], D16[18],
                                            D15[18], D14[18],  D13[18], D12[18], D11[18], D10[18], D9[18],  D8[18],
                                            D7[18],  D6[18],   D5[18],  D4[18],  D3[18],  D2[18],  D1[18],  D0[18]}));
															 
mux_32X1   bit19(.sel(sel), .Y(Y[19]), .D({ D31[19], D30[19],  D29[19], D28[19], D27[19], D26[19], D25[19], D24[19],
                                            D23[19], D22[19],  D21[19], D20[19], D19[19], D18[19], D17[19], D16[19],
                                            D15[19], D14[19],  D13[19], D12[19], D11[19], D10[19], D9[19],  D8[19],
                                            D7[19],  D6[19],   D5[19],  D4[19],  D3[19],  D2[19],  D1[19],  D0[19]}));
															 
mux_32X1   bit20(.sel(sel), .Y(Y[20]), .D({ D31[20], D30[20],  D29[20], D28[20], D27[20], D26[20], D25[20], D24[20],
                                            D23[20], D22[20],  D21[20], D20[20], D19[20], D18[20], D17[20], D16[20],
                                            D15[20], D14[20],  D13[20], D12[20], D11[20], D10[20], D9[20],  D8[20],
                                            D7[20],  D6[20],   D5[20],  D4[20],  D3[20],  D2[20],  D1[20],  D0[20]}));
															 
mux_32X1   bit21(.sel(sel), .Y(Y[21]), .D({ D31[21], D30[21],  D29[21], D28[21], D27[21], D26[21], D25[21], D24[21],
                                            D23[21], D22[21],  D21[21], D20[21], D19[21], D18[21], D17[21], D16[21],
                                            D15[21], D14[21],  D13[21], D12[21], D11[21], D10[21], D9[21],  D8[21],
                                            D7[21],  D6[21],   D5[21],  D4[21],  D3[21],  D2[21],  D1[21],  D0[21]}));
															  
mux_32X1   bit22(.sel(sel), .Y(Y[22]), .D({ D31[22], D30[22],  D29[22], D28[22], D27[22], D26[22], D25[22], D24[22],
                                            D23[22], D22[22],  D21[22], D20[22], D19[22], D18[22], D17[22], D16[22],
                                            D15[22], D14[22],  D13[22], D12[22], D11[22], D10[22], D9[22],  D8[22],
                                            D7[22],  D6[22],   D5[22],  D4[22],  D3[22],  D2[22],  D1[22],  D0[22]}));
															 
mux_32X1   bit23(.sel(sel), .Y(Y[23]), .D({ D31[23], D30[23],  D29[23], D28[23], D27[23], D26[23], D25[23], D24[23],
                                            D23[23], D22[23],  D21[23], D20[23], D19[23], D18[23], D17[23], D16[23],
                                            D15[23], D14[23],  D13[23], D12[23], D11[23], D10[23], D9[23],  D8[23],
                                            D7[23],  D6[23],   D5[23],  D4[23],  D3[23],  D2[23],  D1[23],  D0[23]}));
															 
mux_32X1   bit24(.sel(sel), .Y(Y[24]), .D({ D31[24], D30[24],  D29[24], D28[24], D27[24], D26[24], D25[24], D24[24],
                                            D23[24], D22[24],  D21[24], D20[24], D19[24], D18[24], D17[24], D16[24],
                                            D15[24], D14[24],  D13[24], D12[24], D11[24], D10[24], D9[24],  D8[24],
                                            D7[24],  D6[24],   D5[24],  D4[24],  D3[24],  D2[24],  D1[24],  D0[24]}));
															 
mux_32X1   bit25(.sel(sel), .Y(Y[25]), .D({ D31[25], D30[25],  D29[25], D28[25], D27[25], D26[25], D25[25], D24[25],
                                            D23[25], D22[25],  D21[25], D20[25], D19[25], D18[25], D17[25], D16[25],
                                            D15[25], D14[25],  D13[25], D12[25], D11[25], D10[25], D9[25],  D8[25],
                                            D7[25],  D6[25],   D5[25],  D4[25],  D3[25],  D2[25],  D1[25],  D0[25]}));
															 
mux_32X1   bit26(.sel(sel), .Y(Y[26]), .D({ D31[26], D30[26],  D29[26], D28[26], D27[26], D26[26], D25[26], D24[26],
                                            D23[26], D22[26],  D21[26], D20[26], D19[26], D18[26], D17[26], D16[26],
                                            D15[26], D14[26],  D13[26], D12[26], D11[26], D10[26], D9[26],  D8[26],
                                            D7[26],  D6[26],   D5[26],  D4[26],  D3[26],  D2[26],  D1[26],  D0[26]}));
															 
mux_32X1   bit27(.sel(sel), .Y(Y[27]), .D({ D31[27], D30[27],  D29[27], D28[27], D27[27], D26[27], D25[27], D24[27],
                                            D23[27], D22[27],  D21[27], D20[27], D19[27], D18[27], D17[27], D16[27],
                                            D15[27], D14[27],  D13[27], D12[27], D11[27], D10[27], D9[27],  D8[27],
                                            D7[27],  D6[27],   D5[27],  D4[27],  D3[27],  D2[27],  D1[27],  D0[27]}));
															 
mux_32X1   bit28(.sel(sel), .Y(Y[28]), .D({ D31[28], D30[28],  D29[28], D28[28], D27[28], D26[28], D25[28], D24[28],
                                            D23[28], D22[28],  D21[28], D20[28], D19[28], D18[28], D17[28], D16[28],
                                            D15[28], D14[28],  D13[28], D12[28], D11[28], D10[28], D9[28],  D8[28],
                                            D7[28],  D6[28],   D5[28],  D4[28],  D3[28],  D2[28],  D1[28],  D0[28]}));
															 
mux_32X1   bit29(.sel(sel), .Y(Y[29]), .D({ D31[29], D30[29],  D29[29], D28[29], D27[29], D26[29], D25[29], D24[29],
                                            D23[29], D22[29],  D21[29], D20[29], D19[29], D18[29], D17[29], D16[29],
                                            D15[29], D14[29],  D13[29], D12[29], D11[29], D10[29], D9[29],  D8[29],
                                            D7[29],  D6[29],   D5[29],  D4[29],  D3[29],  D2[29],  D1[29],  D0[29]}));
															 
mux_32X1   bit30(.sel(sel), .Y(Y[30]), .D({ D31[30], D30[30],  D29[30], D28[30], D27[30], D26[30], D25[30], D24[30],
                                            D23[30], D22[30],  D21[30], D20[30], D19[30], D18[30], D17[30], D16[30],
                                            D15[30], D14[30],  D13[30], D12[30], D11[30], D10[30], D9[30],  D8[30],
                                            D7[30],  D6[30],   D5[30],  D4[30],  D3[30],  D2[30],  D1[30],  D0[30]}));
															 
mux_32X1   bit31(.sel(sel), .Y(Y[31]), .D({ D31[31], D30[31],  D29[31], D28[31], D27[31], D26[31], D25[31], D24[31],
                                            D23[31], D22[31],  D21[31], D20[31], D19[31], D18[31], D17[31], D16[31],
                                            D15[31], D14[31],  D13[31], D12[31], D11[31], D10[31], D9[31],  D8[31],
                                            D7[31],  D6[31],   D5[31],  D4[31],  D3[31],  D2[31],  D1[31],  D0[31]}));
															 
endmodule

